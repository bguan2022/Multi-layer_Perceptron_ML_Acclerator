module LUT(
  clk,rst,
  ready,layer2_ready, //ready = layer1_ready
  Input1,Input2,Input3,Input4,Input5,Input6,Input7,Input8,Input9,Input10,Input11,
  Y,Y2,done,Y_sample
);

input clk,rst;
input ready,layer2_ready;
input [15:0] Input1,Input2,Input3,Input4,Input5,Input6,Input7,Input8,Input9,Input10,Input11;
output reg [15:0] Y,Y2;
output reg done;
reg [15:0] X,X2,X3,X4,X5,X6,X7,X8,X9,X10,X11;
//reg [15:0] X,X2;
reg [3:0]cnt;
output reg Y_sample;

// always @(negedge clk ) begin
  // if (rst) begin
    // X<=0;
    // X2<= 0;
    // X3<= 0;
    // X4<= 0;
    // X5<= 0;
    // X6<= 0;
    // X7<= 0;
    // X8<= 0;
    // X9<= 0;
    // X10<= 0;
    // X11<= 0;
  // end else begin
    // if (ready) begin
      // X <= Input1; 
      // if (layer2_ready) begin              
        // X2<= Input2;
        // X3<= Input3;
        // X4<= Input4;
        // X5<= Input5;
        // X6<= Input6;
        // X7<= Input7;
        // X8<= Input8;
        // X9<= Input9;
        // X10<= Input10;
        // X11<= Input11; 
      // end 
	  // else begin
        // X2<= 0;
        // X3<= 0;
        // X4<= 0;
        // X5<= 0;
        // X6<= 0;
        // X7<= 0;
        // X8<= 0;
        // X9<= 0;
        // X10<= 0;
        // X11<= 0;
      // end
    // end else begin
      // X<=X;
      // X2<=X3;
      // X3<=X4;
      // X4<=X5;
      // X5<=X6;
      // X6<=X7;
      // X7<=X8;
      // X8<=X9;
      // X9<=X10;
      // X10<=X11;
      // X11<=0;
    // end
  // end
// end

always @(negedge clk ) begin
  if (rst) begin
    X<=0;
  end 
  else begin
    if (ready) begin
      X <= Input1; 
    end 
	else begin
      X<=X;
    end
  end
end

always @(negedge clk ) begin
  if (rst) begin
    X2<= 0;
    X3<= 0;
    X4<= 0;
    X5<= 0;
    X6<= 0;
    X7<= 0;
    X8<= 0;
    X9<= 0;
    X10<= 0;
    X11<= 0;
  end 
  else begin
    if (layer2_ready && ready) begin
        X2<= Input2;
        X3<= Input3;
        X4<= Input4;
        X5<= Input5;
        X6<= Input6;
        X7<= Input7;
        X8<= Input8;
        X9<= Input9;
        X10<= Input10;
        X11<= Input11;  
    end 
	else begin
      X2<=X3;
      X3<=X4;
      X4<=X5;
      X5<=X6;
      X6<=X7;
      X7<=X8;
      X8<=X9;
      X9<=X10;
      X10<=X11;
      X11<=0;
    end
  end
end





always @(posedge clk) begin
  if (rst) begin
    Y <= 0;
    Y_sample <= 0;
  end else begin
  if (ready) begin
    Y_sample <= 1;
    if (X[15]) begin //negative
      if (X[14:0]<=15'b111101000000000+4'b1101) Y <= 16'b0000000000000000;
      if (X[14:0]>15'b111101000000000+4'b1101 && X[14:0]<=15'b111101000011010+4'b1101) Y <= 16'b0000000000000001;
      if (X[14:0]>15'b111101000011010+4'b1101 && X[14:0]<=15'b111101000110011+4'b1101) Y <= 16'b0000000000000001;
      if (X[14:0]>15'b111101000110011+4'b1101 && X[14:0]<=15'b111101001001101+4'b1101) Y <= 16'b0000000000000001;
      if (X[14:0]>15'b111101001001101+4'b1101 && X[14:0]<=15'b111101001100110+4'b1101) Y <= 16'b0000000000000001;
      if (X[14:0]>15'b111101001100110+4'b1101 && X[14:0]<=15'b111101010000000+4'b1101) Y <= 16'b0000000000000001;
      if (X[14:0]>15'b111101010000000+4'b1101 && X[14:0]<=15'b111101010011010+4'b1101) Y <= 16'b0000000000000001;
      if (X[14:0]>15'b111101010011010+4'b1101 && X[14:0]<=15'b111101010110011+4'b1101) Y <= 16'b0000000000000001;
      if (X[14:0]>15'b111101010110011+4'b1101 && X[14:0]<=15'b111101011001101+4'b1101) Y <= 16'b0000000000000001;
      if (X[14:0]>15'b111101011001101+4'b1101 && X[14:0]<=15'b111101011100110+4'b1101) Y <= 16'b0000000000000010;
      if (X[14:0]>15'b111101011100110+4'b1101 && X[14:0]<=15'b111101100000000+4'b1101) Y <= 16'b0000000000000010;
      if (X[14:0]>15'b111101100000000+4'b1101 && X[14:0]<=15'b111101100011010+4'b1101) Y <= 16'b0000000000000010;
      if (X[14:0]>15'b111101100011010+4'b1101 && X[14:0]<=15'b111101100110011+4'b1101) Y <= 16'b0000000000000010;
      if (X[14:0]>15'b111101100110011+4'b1101 && X[14:0]<=15'b111101101001101+4'b1101) Y <= 16'b0000000000000010;
      if (X[14:0]>15'b111101101001101+4'b1101 && X[14:0]<=15'b111101101100110+4'b1101) Y <= 16'b0000000000000011;
      if (X[14:0]>15'b111101101100110+4'b1101 && X[14:0]<=15'b111101110000000+4'b1101) Y <= 16'b0000000000000011;
      if (X[14:0]>15'b111101110000000+4'b1101 && X[14:0]<=15'b111101110011010+4'b1101) Y <= 16'b0000000000000011;
      if (X[14:0]>15'b111101110011010+4'b1101 && X[14:0]<=15'b111101110110011+4'b1101) Y <= 16'b0000000000000011;
      if (X[14:0]>15'b111101110110011+4'b1101 && X[14:0]<=15'b111101111001101+4'b1101) Y <= 16'b0000000000000100;
      if (X[14:0]>15'b111101111001101+4'b1101 && X[14:0]<=15'b111101111100110+4'b1101) Y <= 16'b0000000000000100;
      if (X[14:0]>15'b111101111100110+4'b1101 && X[14:0]<=15'b111110000000000+4'b1101) Y <= 16'b0000000000000101;
      if (X[14:0]>15'b111110000000000+4'b1101 && X[14:0]<=15'b111110000011010+4'b1101) Y <= 16'b0000000000000101;
      if (X[14:0]>15'b111110000011010+4'b1101 && X[14:0]<=15'b111110000110011+4'b1101) Y <= 16'b0000000000000110;
      if (X[14:0]>15'b111110000110011+4'b1101 && X[14:0]<=15'b111110001001101+4'b1101) Y <= 16'b0000000000000110;
      if (X[14:0]>15'b111110001001101+4'b1101 && X[14:0]<=15'b111110001100110+4'b1101) Y <= 16'b0000000000000111;
      if (X[14:0]>15'b111110001100110+4'b1101 && X[14:0]<=15'b111110010000000+4'b1101) Y <= 16'b0000000000001000;
      if (X[14:0]>15'b111110010000000+4'b1101 && X[14:0]<=15'b111110010011010+4'b1101) Y <= 16'b0000000000001000;
      if (X[14:0]>15'b111110010011010+4'b1101 && X[14:0]<=15'b111110010110011+4'b1101) Y <= 16'b0000000000001001;
      if (X[14:0]>15'b111110010110011+4'b1101 && X[14:0]<=15'b111110011001101+4'b1101) Y <= 16'b0000000000001010;
      if (X[14:0]>15'b111110011001101+4'b1101 && X[14:0]<=15'b111110011100110+4'b1101) Y <= 16'b0000000000001011;
      if (X[14:0]>15'b111110011100110+4'b1101 && X[14:0]<=15'b111110100000000+4'b1101) Y <= 16'b0000000000001100;
      if (X[14:0]>15'b111110100000000+4'b1101 && X[14:0]<=15'b111110100011010+4'b1101) Y <= 16'b0000000000001101;
      if (X[14:0]>15'b111110100011010+4'b1101 && X[14:0]<=15'b111110100110011+4'b1101) Y <= 16'b0000000000001111;
      if (X[14:0]>15'b111110100110011+4'b1101 && X[14:0]<=15'b111110101001101+4'b1101) Y <= 16'b0000000000010000;
      if (X[14:0]>15'b111110101001101+4'b1101 && X[14:0]<=15'b111110101100110+4'b1101) Y <= 16'b0000000000010010;
      if (X[14:0]>15'b111110101100110+4'b1101 && X[14:0]<=15'b111110110000000+4'b1101) Y <= 16'b0000000000010011;
      if (X[14:0]>15'b111110110000000+4'b1101 && X[14:0]<=15'b111110110011010+4'b1101) Y <= 16'b0000000000010101;
      if (X[14:0]>15'b111110110011010+4'b1101 && X[14:0]<=15'b111110110110011+4'b1101) Y <= 16'b0000000000010111;
      if (X[14:0]>15'b111110110110011+4'b1101 && X[14:0]<=15'b111110111001101+4'b1101) Y <= 16'b0000000000011010;
      if (X[14:0]>15'b111110111001101+4'b1101 && X[14:0]<=15'b111110111100110+4'b1101) Y <= 16'b0000000000011100;
      if (X[14:0]>15'b111110111100110+4'b1101 && X[14:0]<=15'b111111000000000+4'b1101) Y <= 16'b0000000000011111;
      if (X[14:0]>15'b111111000000000+4'b1101 && X[14:0]<=15'b111111000011010+4'b1101) Y <= 16'b0000000000100001;
      if (X[14:0]>15'b111111000011010+4'b1101 && X[14:0]<=15'b111111000110011+4'b1101) Y <= 16'b0000000000100100;
      if (X[14:0]>15'b111111000110011+4'b1101 && X[14:0]<=15'b111111001001101+4'b1101) Y <= 16'b0000000000101000;
      if (X[14:0]>15'b111111001001101+4'b1101 && X[14:0]<=15'b111111001100110+4'b1101) Y <= 16'b0000000000101011;
      if (X[14:0]>15'b111111001100110+4'b1101 && X[14:0]<=15'b111111010000000+4'b1101) Y <= 16'b0000000000101111;
      if (X[14:0]>15'b111111010000000+4'b1101 && X[14:0]<=15'b111111010011010+4'b1101) Y <= 16'b0000000000110011;
      if (X[14:0]>15'b111111010011010+4'b1101 && X[14:0]<=15'b111111010110011+4'b1101) Y <= 16'b0000000000110111;
      if (X[14:0]>15'b111111010110011+4'b1101 && X[14:0]<=15'b111111011001101+4'b1101) Y <= 16'b0000000000111011;
      if (X[14:0]>15'b111111011001101+4'b1101 && X[14:0]<=15'b111111011100110+4'b1101) Y <= 16'b0000000001000000;
      if (X[14:0]>15'b111111011100110+4'b1101 && X[14:0]<=15'b111111100000000+4'b1101) Y <= 16'b0000000001000101;
      if (X[14:0]>15'b111111100000000+4'b1101 && X[14:0]<=15'b111111100011010+4'b1101) Y <= 16'b0000000001001010;
      if (X[14:0]>15'b111111100011010+4'b1101 && X[14:0]<=15'b111111100110011+4'b1101) Y <= 16'b0000000001001111;
      if (X[14:0]>15'b111111100110011+4'b1101 && X[14:0]<=15'b111111101001101+4'b1101) Y <= 16'b0000000001010101;
      if (X[14:0]>15'b111111101001101+4'b1101 && X[14:0]<=15'b111111101100110+4'b1101) Y <= 16'b0000000001011011;
      if (X[14:0]>15'b111111101100110+4'b1101 && X[14:0]<=15'b111111110000000+4'b1101) Y <= 16'b0000000001100001;
      if (X[14:0]>15'b111111110000000+4'b1101 && X[14:0]<=15'b111111110011010+4'b1101) Y <= 16'b0000000001100111;
      if (X[14:0]>15'b111111110011010+4'b1101 && X[14:0]<=15'b111111110110011+4'b1101) Y <= 16'b0000000001101101;
      if (X[14:0]>15'b111111110110011+4'b1101 && X[14:0]<=15'b111111111001101+4'b1101) Y <= 16'b0000000001110011;
      if (X[14:0]>15'b111111111001101+4'b1101 && X[14:0]<=15'b111111111100110+4'b1101) Y <= 16'b0000000001111010;
      if (X[14:0]>15'b111111111100110+4'b1101 && X[14:0]<=15'b111111111111111) Y <= 16'b0000000010000000;
    end else begin //positive
      if (X[14:0]>=15'b000011000000000-4'b1101) Y <= 16'b0000000100000000;
      if (X[14:0]>=15'b000000000000000 && X[14:0]<15'b000000000011010-4'b1101) Y <= 16'b0000000010000000;
      if (X[14:0]>=15'b000000000011010-4'b1101 && X[14:0]<15'b000000000110011-4'b1101) Y <= 16'b0000000010000110;
      if (X[14:0]>=15'b000000000110011-4'b1101 && X[14:0]<15'b000000001001101-4'b1101) Y <= 16'b0000000010001101;
      if (X[14:0]>=15'b000000001001101-4'b1101 && X[14:0]<15'b000000001100110-4'b1101) Y <= 16'b0000000010010011;
      if (X[14:0]>=15'b000000001100110-4'b1101 && X[14:0]<15'b000000010000000-4'b1101) Y <= 16'b0000000010011001;
      if (X[14:0]>=15'b000000010000000-4'b1101 && X[14:0]<15'b000000010011010-4'b1101) Y <= 16'b0000000010011111;
      if (X[14:0]>=15'b000000010011010-4'b1101 && X[14:0]<15'b000000010110011-4'b1101) Y <= 16'b0000000010100101;
      if (X[14:0]>=15'b000000010110011-4'b1101 && X[14:0]<15'b000000011001101-4'b1101) Y <= 16'b0000000010101011;
      if (X[14:0]>=15'b000000011001101-4'b1101 && X[14:0]<15'b000000011100110-4'b1101) Y <= 16'b0000000010110001;
      if (X[14:0]>=15'b000000011100110-4'b1101 && X[14:0]<15'b000000100000000-4'b1101) Y <= 16'b0000000010110110;
      if (X[14:0]>=15'b000000100000000-4'b1101 && X[14:0]<15'b000000100011010-4'b1101) Y <= 16'b0000000010111011;
      if (X[14:0]>=15'b000000100011010-4'b1101 && X[14:0]<15'b000000100110011-4'b1101) Y <= 16'b0000000011000000;
      if (X[14:0]>=15'b000000100110011-4'b1101 && X[14:0]<15'b000000101001101-4'b1101) Y <= 16'b0000000011000101;
      if (X[14:0]>=15'b000000101001101-4'b1101 && X[14:0]<15'b000000101100110-4'b1101) Y <= 16'b0000000011001001;
      if (X[14:0]>=15'b000000101100110-4'b1101 && X[14:0]<15'b000000110000000-4'b1101) Y <= 16'b0000000011001101;
      if (X[14:0]>=15'b000000110000000-4'b1101 && X[14:0]<15'b000000110011010-4'b1101) Y <= 16'b0000000011010001;
      if (X[14:0]>=15'b000000110011010-4'b1101 && X[14:0]<15'b000000110110011-4'b1101) Y <= 16'b0000000011010101;
      if (X[14:0]>=15'b000000110110011-4'b1101 && X[14:0]<15'b000000111001101-4'b1101) Y <= 16'b0000000011011000;
      if (X[14:0]>=15'b000000111001101-4'b1101 && X[14:0]<15'b000000111100110-4'b1101) Y <= 16'b0000000011011100;
      if (X[14:0]>=15'b000000111100110-4'b1101 && X[14:0]<15'b000001000000000-4'b1101) Y <= 16'b0000000011011111;
      if (X[14:0]>=15'b000001000000000-4'b1101 && X[14:0]<15'b000001000011010-4'b1101) Y <= 16'b0000000011100001;
      if (X[14:0]>=15'b000001000011010-4'b1101 && X[14:0]<15'b000001000110011-4'b1101) Y <= 16'b0000000011100100;
      if (X[14:0]>=15'b000001000110011-4'b1101 && X[14:0]<15'b000001001001101-4'b1101) Y <= 16'b0000000011100110;
      if (X[14:0]>=15'b000001001001101-4'b1101 && X[14:0]<15'b000001001100110-4'b1101) Y <= 16'b0000000011101001;
      if (X[14:0]>=15'b000001001100110-4'b1101 && X[14:0]<15'b000001010000000-4'b1101) Y <= 16'b0000000011101011;
      if (X[14:0]>=15'b000001010000000-4'b1101 && X[14:0]<15'b000001010011010-4'b1101) Y <= 16'b0000000011101101;
      if (X[14:0]>=15'b000001010011010-4'b1101 && X[14:0]<15'b000001010110011-4'b1101) Y <= 16'b0000000011101110;
      if (X[14:0]>=15'b000001010110011-4'b1101 && X[14:0]<15'b000001011001101-4'b1101) Y <= 16'b0000000011110000;
      if (X[14:0]>=15'b000001011001101-4'b1101 && X[14:0]<15'b000001011100110-4'b1101) Y <= 16'b0000000011110001;
      if (X[14:0]>=15'b000001011100110-4'b1101 && X[14:0]<15'b000001100000000-4'b1101) Y <= 16'b0000000011110011;
      if (X[14:0]>=15'b000001100000000-4'b1101 && X[14:0]<15'b000001100011010-4'b1101) Y <= 16'b0000000011110100;
      if (X[14:0]>=15'b000001100011010-4'b1101 && X[14:0]<15'b000001100110011-4'b1101) Y <= 16'b0000000011110101;
      if (X[14:0]>=15'b000001100110011-4'b1101 && X[14:0]<15'b000001101001101-4'b1101) Y <= 16'b0000000011110110;
      if (X[14:0]>=15'b000001101001101-4'b1101 && X[14:0]<15'b000001101100110-4'b1101) Y <= 16'b0000000011110111;
      if (X[14:0]>=15'b000001101100110-4'b1101 && X[14:0]<15'b000001110000000-4'b1101) Y <= 16'b0000000011111000;
      if (X[14:0]>=15'b000001110000000-4'b1101 && X[14:0]<15'b000001110011010-4'b1101) Y <= 16'b0000000011111000;
      if (X[14:0]>=15'b000001110011010-4'b1101 && X[14:0]<15'b000001110110011-4'b1101) Y <= 16'b0000000011111001;
      if (X[14:0]>=15'b000001110110011-4'b1101 && X[14:0]<15'b000001111001101-4'b1101) Y <= 16'b0000000011111010;
      if (X[14:0]>=15'b000001111001101-4'b1101 && X[14:0]<15'b000001111100110-4'b1101) Y <= 16'b0000000011111010;
      if (X[14:0]>=15'b000001111100110-4'b1101 && X[14:0]<15'b000010000000000-4'b1101) Y <= 16'b0000000011111011;
      if (X[14:0]>=15'b000010000000000-4'b1101 && X[14:0]<15'b000010000011010-4'b1101) Y <= 16'b0000000011111011;
      if (X[14:0]>=15'b000010000011010-4'b1101 && X[14:0]<15'b000010000110011-4'b1101) Y <= 16'b0000000011111100;
      if (X[14:0]>=15'b000010000110011-4'b1101 && X[14:0]<15'b000010001001101-4'b1101) Y <= 16'b0000000011111100;
      if (X[14:0]>=15'b000010001001101-4'b1101 && X[14:0]<15'b000010001100110-4'b1101) Y <= 16'b0000000011111101;
      if (X[14:0]>=15'b000010001100110-4'b1101 && X[14:0]<15'b000010010000000-4'b1101) Y <= 16'b0000000011111101;
      if (X[14:0]>=15'b000010010000000-4'b1101 && X[14:0]<15'b000010010011010-4'b1101) Y <= 16'b0000000011111101;
      if (X[14:0]>=15'b000010010011010-4'b1101 && X[14:0]<15'b000010010110011-4'b1101) Y <= 16'b0000000011111101;
      if (X[14:0]>=15'b000010010110011-4'b1101 && X[14:0]<15'b000010011001101-4'b1101) Y <= 16'b0000000011111110;
      if (X[14:0]>=15'b000010011001101-4'b1101 && X[14:0]<15'b000010011100110-4'b1101) Y <= 16'b0000000011111110;
      if (X[14:0]>=15'b000010011100110-4'b1101 && X[14:0]<15'b000010100000000-4'b1101) Y <= 16'b0000000011111110;
      if (X[14:0]>=15'b000010100000000-4'b1101 && X[14:0]<15'b000010100011010-4'b1101) Y <= 16'b0000000011111110;
      if (X[14:0]>=15'b000010100011010-4'b1101 && X[14:0]<15'b000010100110011-4'b1101) Y <= 16'b0000000011111110;
      if (X[14:0]>=15'b000010100110011-4'b1101 && X[14:0]<15'b000010101001101-4'b1101) Y <= 16'b0000000011111111;
      if (X[14:0]>=15'b000010101001101-4'b1101 && X[14:0]<15'b000010101100110-4'b1101) Y <= 16'b0000000011111111;
      if (X[14:0]>=15'b000010101100110-4'b1101 && X[14:0]<15'b000010110000000-4'b1101) Y <= 16'b0000000011111111;
      if (X[14:0]>=15'b000010110000000-4'b1101 && X[14:0]<15'b000010110011010-4'b1101) Y <= 16'b0000000011111111;
      if (X[14:0]>=15'b000010110011010-4'b1101 && X[14:0]<15'b000010110110011-4'b1101) Y <= 16'b0000000011111111;
      if (X[14:0]>=15'b000010110110011-4'b1101 && X[14:0]<15'b000010111001101-4'b1101) Y <= 16'b0000000011111111;
      if (X[14:0]>=15'b000010111001101-4'b1101 && X[14:0]<15'b000010111100110-4'b1101) Y <= 16'b0000000011111111;
      if (X[14:0]>=15'b000010111100110-4'b1101 && X[14:0]<15'b000011000000000-4'b1101) Y <= 16'b0000000011111111;
    end
  end else begin
    Y <= Y; 
    Y_sample <= 0;
  end
  end
end

always @(posedge clk) begin
  if (rst) begin
    Y2 <= 0;
    done <= 0;
    cnt <= 0;
  end else begin
  if (layer2_ready || (cnt >= 4'd8 && cnt <= 4'd9)) begin
    cnt <= cnt + 1;
    if (X2[15]) begin //negative
      if (X2[14:0]<=15'b111101000000000+4'b1101) Y2 <= 16'b0000000000000000;
      if (X2[14:0]>15'b111101000000000+4'b1101 && X2[14:0]<=15'b111101000011010+4'b1101) Y2 <= 16'b0000000000000001;
      if (X2[14:0]>15'b111101000011010+4'b1101 && X2[14:0]<=15'b111101000110011+4'b1101) Y2 <= 16'b0000000000000001;
      if (X2[14:0]>15'b111101000110011+4'b1101 && X2[14:0]<=15'b111101001001101+4'b1101) Y2 <= 16'b0000000000000001;
      if (X2[14:0]>15'b111101001001101+4'b1101 && X2[14:0]<=15'b111101001100110+4'b1101) Y2 <= 16'b0000000000000001;
      if (X2[14:0]>15'b111101001100110+4'b1101 && X2[14:0]<=15'b111101010000000+4'b1101) Y2 <= 16'b0000000000000001;
      if (X2[14:0]>15'b111101010000000+4'b1101 && X2[14:0]<=15'b111101010011010+4'b1101) Y2 <= 16'b0000000000000001;
      if (X2[14:0]>15'b111101010011010+4'b1101 && X2[14:0]<=15'b111101010110011+4'b1101) Y2 <= 16'b0000000000000001;
      if (X2[14:0]>15'b111101010110011+4'b1101 && X2[14:0]<=15'b111101011001101+4'b1101) Y2 <= 16'b0000000000000001;
      if (X2[14:0]>15'b111101011001101+4'b1101 && X2[14:0]<=15'b111101011100110+4'b1101) Y2 <= 16'b0000000000000010;
      if (X2[14:0]>15'b111101011100110+4'b1101 && X2[14:0]<=15'b111101100000000+4'b1101) Y2 <= 16'b0000000000000010;
      if (X2[14:0]>15'b111101100000000+4'b1101 && X2[14:0]<=15'b111101100011010+4'b1101) Y2 <= 16'b0000000000000010;
      if (X2[14:0]>15'b111101100011010+4'b1101 && X2[14:0]<=15'b111101100110011+4'b1101) Y2 <= 16'b0000000000000010;
      if (X2[14:0]>15'b111101100110011+4'b1101 && X2[14:0]<=15'b111101101001101+4'b1101) Y2 <= 16'b0000000000000010;
      if (X2[14:0]>15'b111101101001101+4'b1101 && X2[14:0]<=15'b111101101100110+4'b1101) Y2 <= 16'b0000000000000011;
      if (X2[14:0]>15'b111101101100110+4'b1101 && X2[14:0]<=15'b111101110000000+4'b1101) Y2 <= 16'b0000000000000011;
      if (X2[14:0]>15'b111101110000000+4'b1101 && X2[14:0]<=15'b111101110011010+4'b1101) Y2 <= 16'b0000000000000011;
      if (X2[14:0]>15'b111101110011010+4'b1101 && X2[14:0]<=15'b111101110110011+4'b1101) Y2 <= 16'b0000000000000011;
      if (X2[14:0]>15'b111101110110011+4'b1101 && X2[14:0]<=15'b111101111001101+4'b1101) Y2 <= 16'b0000000000000100;
      if (X2[14:0]>15'b111101111001101+4'b1101 && X2[14:0]<=15'b111101111100110+4'b1101) Y2 <= 16'b0000000000000100;
      if (X2[14:0]>15'b111101111100110+4'b1101 && X2[14:0]<=15'b111110000000000+4'b1101) Y2 <= 16'b0000000000000101;
      if (X2[14:0]>15'b111110000000000+4'b1101 && X2[14:0]<=15'b111110000011010+4'b1101) Y2 <= 16'b0000000000000101;
      if (X2[14:0]>15'b111110000011010+4'b1101 && X2[14:0]<=15'b111110000110011+4'b1101) Y2 <= 16'b0000000000000110;
      if (X2[14:0]>15'b111110000110011+4'b1101 && X2[14:0]<=15'b111110001001101+4'b1101) Y2 <= 16'b0000000000000110;
      if (X2[14:0]>15'b111110001001101+4'b1101 && X2[14:0]<=15'b111110001100110+4'b1101) Y2 <= 16'b0000000000000111;
      if (X2[14:0]>15'b111110001100110+4'b1101 && X2[14:0]<=15'b111110010000000+4'b1101) Y2 <= 16'b0000000000001000;
      if (X2[14:0]>15'b111110010000000+4'b1101 && X2[14:0]<=15'b111110010011010+4'b1101) Y2 <= 16'b0000000000001000;
      if (X2[14:0]>15'b111110010011010+4'b1101 && X2[14:0]<=15'b111110010110011+4'b1101) Y2 <= 16'b0000000000001001;
      if (X2[14:0]>15'b111110010110011+4'b1101 && X2[14:0]<=15'b111110011001101+4'b1101) Y2 <= 16'b0000000000001010;
      if (X2[14:0]>15'b111110011001101+4'b1101 && X2[14:0]<=15'b111110011100110+4'b1101) Y2 <= 16'b0000000000001011;
      if (X2[14:0]>15'b111110011100110+4'b1101 && X2[14:0]<=15'b111110100000000+4'b1101) Y2 <= 16'b0000000000001100;
      if (X2[14:0]>15'b111110100000000+4'b1101 && X2[14:0]<=15'b111110100011010+4'b1101) Y2 <= 16'b0000000000001101;
      if (X2[14:0]>15'b111110100011010+4'b1101 && X2[14:0]<=15'b111110100110011+4'b1101) Y2 <= 16'b0000000000001111;
      if (X2[14:0]>15'b111110100110011+4'b1101 && X2[14:0]<=15'b111110101001101+4'b1101) Y2 <= 16'b0000000000010000;
      if (X2[14:0]>15'b111110101001101+4'b1101 && X2[14:0]<=15'b111110101100110+4'b1101) Y2 <= 16'b0000000000010010;
      if (X2[14:0]>15'b111110101100110+4'b1101 && X2[14:0]<=15'b111110110000000+4'b1101) Y2 <= 16'b0000000000010011;
      if (X2[14:0]>15'b111110110000000+4'b1101 && X2[14:0]<=15'b111110110011010+4'b1101) Y2 <= 16'b0000000000010101;
      if (X2[14:0]>15'b111110110011010+4'b1101 && X2[14:0]<=15'b111110110110011+4'b1101) Y2 <= 16'b0000000000010111;
      if (X2[14:0]>15'b111110110110011+4'b1101 && X2[14:0]<=15'b111110111001101+4'b1101) Y2 <= 16'b0000000000011010;
      if (X2[14:0]>15'b111110111001101+4'b1101 && X2[14:0]<=15'b111110111100110+4'b1101) Y2 <= 16'b0000000000011100;
      if (X2[14:0]>15'b111110111100110+4'b1101 && X2[14:0]<=15'b111111000000000+4'b1101) Y2 <= 16'b0000000000011111;
      if (X2[14:0]>15'b111111000000000+4'b1101 && X2[14:0]<=15'b111111000011010+4'b1101) Y2 <= 16'b0000000000100001;
      if (X2[14:0]>15'b111111000011010+4'b1101 && X2[14:0]<=15'b111111000110011+4'b1101) Y2 <= 16'b0000000000100100;
      if (X2[14:0]>15'b111111000110011+4'b1101 && X2[14:0]<=15'b111111001001101+4'b1101) Y2 <= 16'b0000000000101000;
      if (X2[14:0]>15'b111111001001101+4'b1101 && X2[14:0]<=15'b111111001100110+4'b1101) Y2 <= 16'b0000000000101011;
      if (X2[14:0]>15'b111111001100110+4'b1101 && X2[14:0]<=15'b111111010000000+4'b1101) Y2 <= 16'b0000000000101111;
      if (X2[14:0]>15'b111111010000000+4'b1101 && X2[14:0]<=15'b111111010011010+4'b1101) Y2 <= 16'b0000000000110011;
      if (X2[14:0]>15'b111111010011010+4'b1101 && X2[14:0]<=15'b111111010110011+4'b1101) Y2 <= 16'b0000000000110111;
      if (X2[14:0]>15'b111111010110011+4'b1101 && X2[14:0]<=15'b111111011001101+4'b1101) Y2 <= 16'b0000000000111011;
      if (X2[14:0]>15'b111111011001101+4'b1101 && X2[14:0]<=15'b111111011100110+4'b1101) Y2 <= 16'b0000000001000000;
      if (X2[14:0]>15'b111111011100110+4'b1101 && X2[14:0]<=15'b111111100000000+4'b1101) Y2 <= 16'b0000000001000101;
      if (X2[14:0]>15'b111111100000000+4'b1101 && X2[14:0]<=15'b111111100011010+4'b1101) Y2 <= 16'b0000000001001010;
      if (X2[14:0]>15'b111111100011010+4'b1101 && X2[14:0]<=15'b111111100110011+4'b1101) Y2 <= 16'b0000000001001111;
      if (X2[14:0]>15'b111111100110011+4'b1101 && X2[14:0]<=15'b111111101001101+4'b1101) Y2 <= 16'b0000000001010101;
      if (X2[14:0]>15'b111111101001101+4'b1101 && X2[14:0]<=15'b111111101100110+4'b1101) Y2 <= 16'b0000000001011011;
      if (X2[14:0]>15'b111111101100110+4'b1101 && X2[14:0]<=15'b111111110000000+4'b1101) Y2 <= 16'b0000000001100001;
      if (X2[14:0]>15'b111111110000000+4'b1101 && X2[14:0]<=15'b111111110011010+4'b1101) Y2 <= 16'b0000000001100111;
      if (X2[14:0]>15'b111111110011010+4'b1101 && X2[14:0]<=15'b111111110110011+4'b1101) Y2 <= 16'b0000000001101101;
      if (X2[14:0]>15'b111111110110011+4'b1101 && X2[14:0]<=15'b111111111001101+4'b1101) Y2 <= 16'b0000000001110011;
      if (X2[14:0]>15'b111111111001101+4'b1101 && X2[14:0]<=15'b111111111100110+4'b1101) Y2 <= 16'b0000000001111010;
      if (X2[14:0]>15'b111111111100110+4'b1101 && X2[14:0]<=15'b111111111111111) Y2 <= 16'b0000000010000000;
    end else begin //positive
      if (X2[14:0]>=15'b000011000000000-4'b1101) Y2 <= 16'b0000000100000000;
      if (X2[14:0]>=15'b000000000000000 && X2[14:0]<15'b000000000011010-4'b1101) Y2 <= 16'b0000000010000000;
      if (X2[14:0]>=15'b000000000011010-4'b1101 && X2[14:0]<15'b000000000110011-4'b1101) Y2 <= 16'b0000000010000110;
      if (X2[14:0]>=15'b000000000110011-4'b1101 && X2[14:0]<15'b000000001001101-4'b1101) Y2 <= 16'b0000000010001101;
      if (X2[14:0]>=15'b000000001001101-4'b1101 && X2[14:0]<15'b000000001100110-4'b1101) Y2 <= 16'b0000000010010011;
      if (X2[14:0]>=15'b000000001100110-4'b1101 && X2[14:0]<15'b000000010000000-4'b1101) Y2 <= 16'b0000000010011001;
      if (X2[14:0]>=15'b000000010000000-4'b1101 && X2[14:0]<15'b000000010011010-4'b1101) Y2 <= 16'b0000000010011111;
      if (X2[14:0]>=15'b000000010011010-4'b1101 && X2[14:0]<15'b000000010110011-4'b1101) Y2 <= 16'b0000000010100101;
      if (X2[14:0]>=15'b000000010110011-4'b1101 && X2[14:0]<15'b000000011001101-4'b1101) Y2 <= 16'b0000000010101011;
      if (X2[14:0]>=15'b000000011001101-4'b1101 && X2[14:0]<15'b000000011100110-4'b1101) Y2 <= 16'b0000000010110001;
      if (X2[14:0]>=15'b000000011100110-4'b1101 && X2[14:0]<15'b000000100000000-4'b1101) Y2 <= 16'b0000000010110110;
      if (X2[14:0]>=15'b000000100000000-4'b1101 && X2[14:0]<15'b000000100011010-4'b1101) Y2 <= 16'b0000000010111011;
      if (X2[14:0]>=15'b000000100011010-4'b1101 && X2[14:0]<15'b000000100110011-4'b1101) Y2 <= 16'b0000000011000000;
      if (X2[14:0]>=15'b000000100110011-4'b1101 && X2[14:0]<15'b000000101001101-4'b1101) Y2 <= 16'b0000000011000101;
      if (X2[14:0]>=15'b000000101001101-4'b1101 && X2[14:0]<15'b000000101100110-4'b1101) Y2 <= 16'b0000000011001001;
      if (X2[14:0]>=15'b000000101100110-4'b1101 && X2[14:0]<15'b000000110000000-4'b1101) Y2 <= 16'b0000000011001101;
      if (X2[14:0]>=15'b000000110000000-4'b1101 && X2[14:0]<15'b000000110011010-4'b1101) Y2 <= 16'b0000000011010001;
      if (X2[14:0]>=15'b000000110011010-4'b1101 && X2[14:0]<15'b000000110110011-4'b1101) Y2 <= 16'b0000000011010101;
      if (X2[14:0]>=15'b000000110110011-4'b1101 && X2[14:0]<15'b000000111001101-4'b1101) Y2 <= 16'b0000000011011000;
      if (X2[14:0]>=15'b000000111001101-4'b1101 && X2[14:0]<15'b000000111100110-4'b1101) Y2 <= 16'b0000000011011100;
      if (X2[14:0]>=15'b000000111100110-4'b1101 && X2[14:0]<15'b000001000000000-4'b1101) Y2 <= 16'b0000000011011111;
      if (X2[14:0]>=15'b000001000000000-4'b1101 && X2[14:0]<15'b000001000011010-4'b1101) Y2 <= 16'b0000000011100001;
      if (X2[14:0]>=15'b000001000011010-4'b1101 && X2[14:0]<15'b000001000110011-4'b1101) Y2 <= 16'b0000000011100100;
      if (X2[14:0]>=15'b000001000110011-4'b1101 && X2[14:0]<15'b000001001001101-4'b1101) Y2 <= 16'b0000000011100110;
      if (X2[14:0]>=15'b000001001001101-4'b1101 && X2[14:0]<15'b000001001100110-4'b1101) Y2 <= 16'b0000000011101001;
      if (X2[14:0]>=15'b000001001100110-4'b1101 && X2[14:0]<15'b000001010000000-4'b1101) Y2 <= 16'b0000000011101011;
      if (X2[14:0]>=15'b000001010000000-4'b1101 && X2[14:0]<15'b000001010011010-4'b1101) Y2 <= 16'b0000000011101101;
      if (X2[14:0]>=15'b000001010011010-4'b1101 && X2[14:0]<15'b000001010110011-4'b1101) Y2 <= 16'b0000000011101110;
      if (X2[14:0]>=15'b000001010110011-4'b1101 && X2[14:0]<15'b000001011001101-4'b1101) Y2 <= 16'b0000000011110000;
      if (X2[14:0]>=15'b000001011001101-4'b1101 && X2[14:0]<15'b000001011100110-4'b1101) Y2 <= 16'b0000000011110001;
      if (X2[14:0]>=15'b000001011100110-4'b1101 && X2[14:0]<15'b000001100000000-4'b1101) Y2 <= 16'b0000000011110011;
      if (X2[14:0]>=15'b000001100000000-4'b1101 && X2[14:0]<15'b000001100011010-4'b1101) Y2 <= 16'b0000000011110100;
      if (X2[14:0]>=15'b000001100011010-4'b1101 && X2[14:0]<15'b000001100110011-4'b1101) Y2 <= 16'b0000000011110101;
      if (X2[14:0]>=15'b000001100110011-4'b1101 && X2[14:0]<15'b000001101001101-4'b1101) Y2 <= 16'b0000000011110110;
      if (X2[14:0]>=15'b000001101001101-4'b1101 && X2[14:0]<15'b000001101100110-4'b1101) Y2 <= 16'b0000000011110111;
      if (X2[14:0]>=15'b000001101100110-4'b1101 && X2[14:0]<15'b000001110000000-4'b1101) Y2 <= 16'b0000000011111000;
      if (X2[14:0]>=15'b000001110000000-4'b1101 && X2[14:0]<15'b000001110011010-4'b1101) Y2 <= 16'b0000000011111000;
      if (X2[14:0]>=15'b000001110011010-4'b1101 && X2[14:0]<15'b000001110110011-4'b1101) Y2 <= 16'b0000000011111001;
      if (X2[14:0]>=15'b000001110110011-4'b1101 && X2[14:0]<15'b000001111001101-4'b1101) Y2 <= 16'b0000000011111010;
      if (X2[14:0]>=15'b000001111001101-4'b1101 && X2[14:0]<15'b000001111100110-4'b1101) Y2 <= 16'b0000000011111010;
      if (X2[14:0]>=15'b000001111100110-4'b1101 && X2[14:0]<15'b000010000000000-4'b1101) Y2 <= 16'b0000000011111011;
      if (X2[14:0]>=15'b000010000000000-4'b1101 && X2[14:0]<15'b000010000011010-4'b1101) Y2 <= 16'b0000000011111011;
      if (X2[14:0]>=15'b000010000011010-4'b1101 && X2[14:0]<15'b000010000110011-4'b1101) Y2 <= 16'b0000000011111100;
      if (X2[14:0]>=15'b000010000110011-4'b1101 && X2[14:0]<15'b000010001001101-4'b1101) Y2 <= 16'b0000000011111100;
      if (X2[14:0]>=15'b000010001001101-4'b1101 && X2[14:0]<15'b000010001100110-4'b1101) Y2 <= 16'b0000000011111101;
      if (X2[14:0]>=15'b000010001100110-4'b1101 && X2[14:0]<15'b000010010000000-4'b1101) Y2 <= 16'b0000000011111101;
      if (X2[14:0]>=15'b000010010000000-4'b1101 && X2[14:0]<15'b000010010011010-4'b1101) Y2 <= 16'b0000000011111101;
      if (X2[14:0]>=15'b000010010011010-4'b1101 && X2[14:0]<15'b000010010110011-4'b1101) Y2 <= 16'b0000000011111101;
      if (X2[14:0]>=15'b000010010110011-4'b1101 && X2[14:0]<15'b000010011001101-4'b1101) Y2 <= 16'b0000000011111110;
      if (X2[14:0]>=15'b000010011001101-4'b1101 && X2[14:0]<15'b000010011100110-4'b1101) Y2 <= 16'b0000000011111110;
      if (X2[14:0]>=15'b000010011100110-4'b1101 && X2[14:0]<15'b000010100000000-4'b1101) Y2 <= 16'b0000000011111110;
      if (X2[14:0]>=15'b000010100000000-4'b1101 && X2[14:0]<15'b000010100011010-4'b1101) Y2 <= 16'b0000000011111110;
      if (X2[14:0]>=15'b000010100011010-4'b1101 && X2[14:0]<15'b000010100110011-4'b1101) Y2 <= 16'b0000000011111110;
      if (X2[14:0]>=15'b000010100110011-4'b1101 && X2[14:0]<15'b000010101001101-4'b1101) Y2 <= 16'b0000000011111111;
      if (X2[14:0]>=15'b000010101001101-4'b1101 && X2[14:0]<15'b000010101100110-4'b1101) Y2 <= 16'b0000000011111111;
      if (X2[14:0]>=15'b000010101100110-4'b1101 && X2[14:0]<15'b000010110000000-4'b1101) Y2 <= 16'b0000000011111111;
      if (X2[14:0]>=15'b000010110000000-4'b1101 && X2[14:0]<15'b000010110011010-4'b1101) Y2 <= 16'b0000000011111111;
      if (X2[14:0]>=15'b000010110011010-4'b1101 && X2[14:0]<15'b000010110110011-4'b1101) Y2 <= 16'b0000000011111111;
      if (X2[14:0]>=15'b000010110110011-4'b1101 && X2[14:0]<15'b000010111001101-4'b1101) Y2 <= 16'b0000000011111111;
      if (X2[14:0]>=15'b000010111001101-4'b1101 && X2[14:0]<15'b000010111100110-4'b1101) Y2 <= 16'b0000000011111111;
      if (X2[14:0]>=15'b000010111100110-4'b1101 && X2[14:0]<15'b000011000000000-4'b1101) Y2 <= 16'b0000000011111111;
    end
    if (cnt<=9) done <= 1;
    else done<=0;
  end else begin
    Y2 <= 0;
    done <= 0;
    cnt <= 0;
  end
  end
end

endmodule // LUT